--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package autoinit_definitions is

 constant scrodpre_len : integer :=3;
 type scrodpre is array (0 to scrodpre_len-1) of std_logic_vector(23 downto 0);
 constant init_scrodpre : scrodpre:= (x"050080",x"060140",x"000000");
 	constant TRIGGER_SCALER_BIT_WIDTH      : integer := 32;

 	constant INIT_CNT1_MAX: integer:=1000000;
	constant WAIT_CNT1_MAX: integer:=1000000;-- wait between regs this long 

  constant scrodpost_len : integer :=35;
  type scrodpost is array (0 to scrodpost_len-1) of std_logic_vector(23 downto 0);
 constant init_scrodpost : scrodpost:= (
 x"140000",
 x"1E0000",
 x"1F0000",
 x"320000",
 x"2C0000",
 x"2D0001",
 x"2D0000",
 x"3301E7",
 x"340000",
 x"350000",
 x"3600A0",	-- digitization window offset (aka look back- LKBK)
 x"370001",
 x"370000",
 x"380000",
 x"390004",
 x"3A0000",
 x"4801E7",
 x"3D0F00",
 x"260000",
 x"260800",
 x"260000",
 x"2610A0",
 x"270000",
 x"0B8001",
 x"0A0000",
 x"0A0001",
 x"0A0000",
 x"3E0000",
 x"460000",
 x"470000",
 x"470001",
 x"470000",
 x"460001",
 x"27C1E7",-- Mask DCs that are not connected
 x"007FFF"
 );

  constant scrodpeds_len : integer :=33;
  type scrodpeds is array (0 to scrodpeds_len-1) of std_logic_vector(23 downto 0);
 constant init_scrodpeds : scrodpeds:= (
 x"140000",
 x"1E0000",
 x"320000",
 x"2C0000",
 x"2D0001",
 x"2D0000",
 x"3303FF",
 x"340000",
 x"350000",
 x"360000",	
 x"370001",
 x"370000",
 x"380000",
 x"390004",
 x"3A0000",
 x"4803FF",
 x"3D0F00",
 x"260000",
 x"260800",
 x"260000",

 x"0B8001",
 x"0A0000",
 x"0A0001",
 x"0A0000",

 x"260000",
 x"264000",
 x"26C000",
 x"264000",
 x"270000",

 x"2AFE00",
 x"2903FF",
 x"2983FF",
 x"2903FF"
 );


 constant asic_trig_threshold:std_logic_vector(15 downto 0):=x"0BB8"; --is 3000 decimal

 constant asicregs_len : integer :=63;
	type asicregs is array (0 to asicregs_len-1) of std_logic_vector(23 downto 0);
 constant init_asicregs : asicregs:=(
 x"00" & asic_trig_threshold,
 x"02" & asic_trig_threshold,
 x"04" & asic_trig_threshold,
 x"06" & asic_trig_threshold,
 x"08" & asic_trig_threshold,
 x"0A" & asic_trig_threshold,
 x"0C" & asic_trig_threshold,
 x"0E" & asic_trig_threshold,
 x"10" & asic_trig_threshold,
 x"12" & asic_trig_threshold,
 x"14" & asic_trig_threshold,
 x"16" & asic_trig_threshold,
 x"18" & asic_trig_threshold,
 x"1A" & asic_trig_threshold,
 x"1C" & asic_trig_threshold,
 x"1E" & asic_trig_threshold,
 x"01" & x"03D9",
 x"03" & x"03D9",
 x"05" & x"03D9",
 x"07" & x"03D9",
 x"09" & x"03D9",
 x"0B" & x"03D9",
 x"0D" & x"03D9",
 x"0F" & x"03D9",
 x"11" & x"03D9",
 x"13" & x"03D9",
 x"15" & x"03D9",
 x"17" & x"03D9",
 x"19" & x"03D9",
 x"1B" & x"03D9",
 x"1D" & x"03D9",
 x"1F" & x"03D9",

 x"30" & x"0514",
 x"31" & x"0000",
 x"32" & x"0A5A",
 x"33" & x"044C",
 x"34" & x"05DC",
 x"35" & x"0426",
 x"36" & x"04B9",
 x"37" & x"0000",
 x"38" & x"0480",
 x"39" & x"0000",
 x"3A" & x"08BB",
 x"3B" & x"0000",
 x"3D" & x"04A6",
 x"3E" & x"044C",
 x"3F" & x"044C",
 x"40" & x"008F",
 x"41" & x"00A3",
 x"42" & x"000D",
 x"43" & x"0021",
 x"44" & x"0014",
 x"45" & x"0028",
 x"46" & x"0021",
 x"47" & x"0035",
 x"48" & x"0038",
 x"49" & x"000C",
 x"4A" & x"0028",
 x"4B" & x"003A",
 x"4C" & x"02E1",
 x"4D" & x"0C28",
 x"4E" & x"0480",
 x"4F" & x"0AAA"

 );
 

constant scrod_rcl_autoinit_len: integer:=1250;
 
type scrod_rcl_autoinit is array (0 to scrod_rcl_autoinit_len-1) of std_logic_vector(31 downto 0);
constant init_scrod_rcl_autoinit : scrod_rcl_autoinit:=(
x"01234567",x"AE000100",x"AF000000",x"AE000100",x"AF008000",x"AE000100",x"AE008000",x"AE000100",
x"AE000100",x"AF00FFFF",x"AE000100",x"AE000100",x"AF008000",x"AE000100",x"AF050080",x"AE000100",
x"AF060140",x"AE000100",x"B00005AA",x"B00205AA",x"B00405AA",x"B00605AA",x"B00805AA",x"B00A05AA",
x"B00C05AA",x"B00E05AA",x"B01005AA",x"B01205AA",x"B01405AA",x"B01605AA",x"B01805AA",x"B01A05AA",
x"B01C05AA",x"B01E05AA",x"B00103D9",x"B00303D9",x"B00503D9",x"B00703D9",x"B00903D9",x"B00B03D9",
x"B00D03D9",x"B00F03D9",x"B01103D9",x"B01303D9",x"B01503D9",x"B01703D9",x"B01903D9",x"B01B03D9",
x"B01D03D9",x"B01F03D9",x"B0300514",x"B0310000",x"B0320A5A",x"B033044C",x"B03405DC",x"B0350426",
x"B03604B9",x"B0370000",x"B0380480",x"B0390000",x"B03A08BB",x"B03B0000",x"B03D04A6",x"B03E044C",
x"B03F044C",x"B040008F",x"B04100A3",x"B042000D",x"B0430021",x"B0440014",x"B0450028",x"B0460021",
x"B0470035",x"B0480038",x"B049000C",x"B04A0028",x"B04B003A",x"B04C02E1",x"B04D0C28",x"B04E0480",
x"B04F0AAA",x"B10005AA",x"B10205AA",x"B10405AA",x"B10605AA",x"B10805AA",x"B10A05AA",x"B10C05AA",
x"B10E05AA",x"B11005AA",x"B11205AA",x"B11405AA",x"B11605AA",x"B11805AA",x"B11A05AA",x"B11C05AA",
x"B11E05AA",x"B10103D9",x"B10303D9",x"B10503D9",x"B10703D9",x"B10903D9",x"B10B03D9",x"B10D03D9",
x"B10F03D9",x"B11103D9",x"B11303D9",x"B11503D9",x"B11703D9",x"B11903D9",x"B11B03D9",x"B11D03D9",
x"B11F03D9",x"B1300514",x"B1310000",x"B1320A5A",x"B133044C",x"B13405DC",x"B1350426",x"B13604B9",
x"B1370000",x"B1380480",x"B1390000",x"B13A08BB",x"B13B0000",x"B13D04A6",x"B13E044C",x"B13F044C",
x"B140008F",x"B14100A3",x"B142000D",x"B1430021",x"B1440014",x"B1450028",x"B1460021",x"B1470035",
x"B1480038",x"B149000C",x"B14A0028",x"B14B003A",x"B14C02E1",x"B14D0C28",x"B14E0480",x"B14F0AAA",
x"B20005AA",x"B20205AA",x"B20405AA",x"B20605AA",x"B20805AA",x"B20A05AA",x"B20C05AA",x"B20E05AA",
x"B21005AA",x"B21205AA",x"B21405AA",x"B21605AA",x"B21805AA",x"B21A05AA",x"B21C05AA",x"B21E05AA",
x"B20103D9",x"B20303D9",x"B20503D9",x"B20703D9",x"B20903D9",x"B20B03D9",x"B20D03D9",x"B20F03D9",
x"B21103D9",x"B21303D9",x"B21503D9",x"B21703D9",x"B21903D9",x"B21B03D9",x"B21D03D9",x"B21F03D9",
x"B2300514",x"B2310000",x"B2320A5A",x"B233044C",x"B23405DC",x"B2350426",x"B23604B9",x"B2370000",
x"B2380480",x"B2390000",x"B23A08BB",x"B23B0000",x"B23D04A6",x"B23E044C",x"B23F044C",x"B240008F",
x"B24100A3",x"B242000D",x"B2430021",x"B2440014",x"B2450028",x"B2460021",x"B2470035",x"B2480038",
x"B249000C",x"B24A0028",x"B24B003A",x"B24C02E1",x"B24D0C28",x"B24E0480",x"B24F0AAA",x"B30005AA",
x"B30205AA",x"B30405AA",x"B30605AA",x"B30805AA",x"B30A05AA",x"B30C05AA",x"B30E05AA",x"B31005AA",
x"B31205AA",x"B31405AA",x"B31605AA",x"B31805AA",x"B31A05AA",x"B31C05AA",x"B31E05AA",x"B30103D9",
x"B30303D9",x"B30503D9",x"B30703D9",x"B30903D9",x"B30B03D9",x"B30D03D9",x"B30F03D9",x"B31103D9",
x"B31303D9",x"B31503D9",x"B31703D9",x"B31903D9",x"B31B03D9",x"B31D03D9",x"B31F03D9",x"B3300514",
x"B3310000",x"B3320A5A",x"B333044C",x"B33405DC",x"B3350426",x"B33604B9",x"B3370000",x"B3380480",
x"B3390000",x"B33A08BB",x"B33B0000",x"B33D04A6",x"B33E044C",x"B33F044C",x"B340008F",x"B34100A3",
x"B342000D",x"B3430021",x"B3440014",x"B3450028",x"B3460021",x"B3470035",x"B3480038",x"B349000C",
x"B34A0028",x"B34B003A",x"B34C02E1",x"B34D0C28",x"B34E0480",x"B34F0AAA",x"B40005AA",x"B40205AA",
x"B40405AA",x"B40605AA",x"B40805AA",x"B40A05AA",x"B40C05AA",x"B40E05AA",x"B41005AA",x"B41205AA",
x"B41405AA",x"B41605AA",x"B41805AA",x"B41A05AA",x"B41C05AA",x"B41E05AA",x"B40103D9",x"B40303D9",
x"B40503D9",x"B40703D9",x"B40903D9",x"B40B03D9",x"B40D03D9",x"B40F03D9",x"B41103D9",x"B41303D9",
x"B41503D9",x"B41703D9",x"B41903D9",x"B41B03D9",x"B41D03D9",x"B41F03D9",x"B4300514",x"B4310000",
x"B4320A5A",x"B433044C",x"B43405DC",x"B4350426",x"B43604B9",x"B4370000",x"B4380480",x"B4390000",
x"B43A08BB",x"B43B0000",x"B43D04A6",x"B43E044C",x"B43F044C",x"B440008F",x"B44100A3",x"B442000D",
x"B4430021",x"B4440014",x"B4450028",x"B4460021",x"B4470035",x"B4480038",x"B449000C",x"B44A0028",
x"B44B003A",x"B44C02E1",x"B44D0C28",x"B44E0480",x"B44F0AAA",x"B50005AA",x"B50205AA",x"B50405AA",
x"B50605AA",x"B50805AA",x"B50A05AA",x"B50C05AA",x"B50E05AA",x"B51005AA",x"B51205AA",x"B51405AA",
x"B51605AA",x"B51805AA",x"B51A05AA",x"B51C05AA",x"B51E05AA",x"B50103D9",x"B50303D9",x"B50503D9",
x"B50703D9",x"B50903D9",x"B50B03D9",x"B50D03D9",x"B50F03D9",x"B51103D9",x"B51303D9",x"B51503D9",
x"B51703D9",x"B51903D9",x"B51B03D9",x"B51D03D9",x"B51F03D9",x"B5300514",x"B5310000",x"B5320A5A",
x"B533044C",x"B53405DC",x"B5350426",x"B53604B9",x"B5370000",x"B5380480",x"B5390000",x"B53A08BB",
x"B53B0000",x"B53D04A6",x"B53E044C",x"B53F044C",x"B540008F",x"B54100A3",x"B542000D",x"B5430021",
x"B5440014",x"B5450028",x"B5460021",x"B5470035",x"B5480038",x"B549000C",x"B54A0028",x"B54B003A",
x"B54C02E1",x"B54D0C28",x"B54E0480",x"B54F0AAA",x"B60005AA",x"B60205AA",x"B60405AA",x"B60605AA",
x"B60805AA",x"B60A05AA",x"B60C05AA",x"B60E05AA",x"B61005AA",x"B61205AA",x"B61405AA",x"B61605AA",
x"B61805AA",x"B61A05AA",x"B61C05AA",x"B61E05AA",x"B60103D9",x"B60303D9",x"B60503D9",x"B60703D9",
x"B60903D9",x"B60B03D9",x"B60D03D9",x"B60F03D9",x"B61103D9",x"B61303D9",x"B61503D9",x"B61703D9",
x"B61903D9",x"B61B03D9",x"B61D03D9",x"B61F03D9",x"B6300514",x"B6310000",x"B6320A5A",x"B633044C",
x"B63405DC",x"B6350426",x"B63604B9",x"B6370000",x"B6380480",x"B6390000",x"B63A08BB",x"B63B0000",
x"B63D04A6",x"B63E044C",x"B63F044C",x"B640008F",x"B64100A3",x"B642000D",x"B6430021",x"B6440014",
x"B6450028",x"B6460021",x"B6470035",x"B6480038",x"B649000C",x"B64A0028",x"B64B003A",x"B64C02E1",
x"B64D0C28",x"B64E0480",x"B64F0AAA",x"B70005AA",x"B70205AA",x"B70405AA",x"B70605AA",x"B70805AA",
x"B70A05AA",x"B70C05AA",x"B70E05AA",x"B71005AA",x"B71205AA",x"B71405AA",x"B71605AA",x"B71805AA",
x"B71A05AA",x"B71C05AA",x"B71E05AA",x"B70103D9",x"B70303D9",x"B70503D9",x"B70703D9",x"B70903D9",
x"B70B03D9",x"B70D03D9",x"B70F03D9",x"B71103D9",x"B71303D9",x"B71503D9",x"B71703D9",x"B71903D9",
x"B71B03D9",x"B71D03D9",x"B71F03D9",x"B7300514",x"B7310000",x"B7320A5A",x"B733044C",x"B73405DC",
x"B7350426",x"B73604B9",x"B7370000",x"B7380480",x"B7390000",x"B73A08BB",x"B73B0000",x"B73D04A6",
x"B73E044C",x"B73F044C",x"B740008F",x"B74100A3",x"B742000D",x"B7430021",x"B7440014",x"B7450028",
x"B7460021",x"B7470035",x"B7480038",x"B749000C",x"B74A0028",x"B74B003A",x"B74C02E1",x"B74D0C28",
x"B74E0480",x"B74F0AAA",x"B80005AA",x"B80205AA",x"B80405AA",x"B80605AA",x"B80805AA",x"B80A05AA",
x"B80C05AA",x"B80E05AA",x"B81005AA",x"B81205AA",x"B81405AA",x"B81605AA",x"B81805AA",x"B81A05AA",
x"B81C05AA",x"B81E05AA",x"B80103D9",x"B80303D9",x"B80503D9",x"B80703D9",x"B80903D9",x"B80B03D9",
x"B80D03D9",x"B80F03D9",x"B81103D9",x"B81303D9",x"B81503D9",x"B81703D9",x"B81903D9",x"B81B03D9",
x"B81D03D9",x"B81F03D9",x"B8300514",x"B8310000",x"B8320A5A",x"B833044C",x"B83405DC",x"B8350426",
x"B83604B9",x"B8370000",x"B8380480",x"B8390000",x"B83A08BB",x"B83B0000",x"B83D04A6",x"B83E044C",
x"B83F044C",x"B840008F",x"B84100A3",x"B842000D",x"B8430021",x"B8440014",x"B8450028",x"B8460021",
x"B8470035",x"B8480038",x"B849000C",x"B84A0028",x"B84B003A",x"B84C02E1",x"B84D0C28",x"B84E0480",
x"B84F0AAA",x"B90005AA",x"B90205AA",x"B90405AA",x"B90605AA",x"B90805AA",x"B90A05AA",x"B90C05AA",
x"B90E05AA",x"B91005AA",x"B91205AA",x"B91405AA",x"B91605AA",x"B91805AA",x"B91A05AA",x"B91C05AA",
x"B91E05AA",x"B90103D9",x"B90303D9",x"B90503D9",x"B90703D9",x"B90903D9",x"B90B03D9",x"B90D03D9",
x"B90F03D9",x"B91103D9",x"B91303D9",x"B91503D9",x"B91703D9",x"B91903D9",x"B91B03D9",x"B91D03D9",
x"B91F03D9",x"B9300514",x"B9310000",x"B9320A5A",x"B933044C",x"B93405DC",x"B9350426",x"B93604B9",
x"B9370000",x"B9380480",x"B9390000",x"B93A08BB",x"B93B0000",x"B93D04A6",x"B93E044C",x"B93F044C",
x"B940008F",x"B94100A3",x"B942000D",x"B9430021",x"B9440014",x"B9450028",x"B9460021",x"B9470035",
x"B9480038",x"B949000C",x"B94A0028",x"B94B003A",x"B94C02E1",x"B94D0C28",x"B94E0480",x"B94F0AAA",
x"C00000FF",x"C00100FF",x"C00200FF",x"C00300FF",x"C00400FF",x"C00500FF",x"C00600FF",x"C00700FF",
x"C00800FF",x"C00900FF",x"C00A00FF",x"C00B00FF",x"C00C00FF",x"C00D00FF",x"C00E00FF",x"C00F00FF",
x"C01000FF",x"C01100FF",x"C01200FF",x"C01300FF",x"C01400FF",x"C01500FF",x"C01600FF",x"C01700FF",
x"C01800FF",x"C01900FF",x"C01A00FF",x"C01B00FF",x"C01C00FF",x"C01D00FF",x"C01E00FF",x"C01F00FF",
x"C02000FF",x"C02100FF",x"C02200FF",x"C02300FF",x"C02400FF",x"C02500FF",x"C02600FF",x"C02700FF",
x"C02800FF",x"C02900FF",x"C02A00FF",x"C02B00FF",x"C02C00FF",x"C02D00FF",x"C02E00FF",x"C02F00FF",
x"C03000FF",x"C03100FF",x"C03200FF",x"C03300FF",x"C03400FF",x"C03500FF",x"C03600FF",x"C03700FF",
x"C03800FF",x"C03900FF",x"C03A00FF",x"C03B00FF",x"C03C00FF",x"C03D00FF",x"C03E00FF",x"C03F00FF",
x"C04000FF",x"C04100FF",x"C04200FF",x"C04300FF",x"C04400FF",x"C04500FF",x"C04600FF",x"C04700FF",
x"C04800FF",x"C04900FF",x"C04A00FF",x"C04B00FF",x"C04C00FF",x"C04D00FF",x"C04E00FF",x"C04F00FF",
x"C05000FF",x"C05100FF",x"C05200FF",x"C05300FF",x"C05400FF",x"C05500FF",x"C05600FF",x"C05700FF",
x"C05800FF",x"C05900FF",x"C05A00FF",x"C05B00FF",x"C05C00FF",x"C05D00FF",x"C05E00FF",x"C05F00FF",
x"C06000FF",x"C06100FF",x"C06200FF",x"C06300FF",x"C06400FF",x"C06500FF",x"C06600FF",x"C06700FF",
x"C06800FF",x"C06900FF",x"C06A00FF",x"C06B00FF",x"C06C00FF",x"C06D00FF",x"C06E00FF",x"C06F00FF",
x"C07000FF",x"C07100FF",x"C07200FF",x"C07300FF",x"C07400FF",x"C07500FF",x"C07600FF",x"C07700FF",
x"C07800FF",x"C07900FF",x"C07A00FF",x"C07B00FF",x"C07C00FF",x"C07D00FF",x"C07E00FF",x"C07F00FF",
x"C08000FF",x"C08100FF",x"C08200FF",x"C08300FF",x"C08400FF",x"C08500FF",x"C08600FF",x"C08700FF",
x"C08800FF",x"C08900FF",x"C08A00FF",x"C08B00FF",x"C08C00FF",x"C08D00FF",x"C08E00FF",x"C08F00FF",
x"C09000FF",x"C09100FF",x"C09200FF",x"C09300FF",x"C09400FF",x"C09500FF",x"C09600FF",x"C09700FF",
x"C09800FF",x"C09900FF",x"C09A00FF",x"C09B00FF",x"C09C00FF",x"C09D00FF",x"C09E00FF",x"C09F00FF",
x"AF4D0000",x"AE000100",x"AF140000",x"AE000100",x"AF1E0000",x"AE000100",x"AF320000",x"AE000100",
x"AF2C0000",x"AE000100",x"AF2D0001",x"AE000100",x"AF2D0000",x"AE000100",x"AF3303FF",x"AE000100",
x"AF340000",x"AE000100",x"AF350000",x"AE000100",x"AF360000",x"AE000100",x"AF370001",x"AE000100",
x"AF370000",x"AE000100",x"AF380000",x"AE000100",x"AF390004",x"AE000100",x"AF3A0000",x"AE000100",
x"AF4803FF",x"AE000100",x"AF3D0F00",x"AE000100",x"AF260000",x"AE000100",x"AF260800",x"AE000100",
x"AF260000",x"AE000100",x"AF0B8001",x"AE000100",x"AF0A0000",x"AE000100",x"AF0A0001",x"AE000100",
x"AF0A0000",x"AE000100",x"AF260000",x"AE000100",x"AF264000",x"AE000100",x"AF26C000",x"AE000100",
x"AF264000",x"AE000100",x"AF270000",x"AE000100",x"AF2AFE00",x"AE000100",x"AF290200",x"AE000100",
x"AF298200",x"AE00FFFF",x"AF290200",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",
x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AF4D0000",x"AE000100",x"AF140000",x"AE000100",
x"AF1E0000",x"AE000100",x"AF320000",x"AE000100",x"AF2C0000",x"AE000100",x"AF2D0001",x"AE000100",
x"AF2D0000",x"AE000100",x"AF3303FF",x"AE000100",x"AF340000",x"AE000100",x"AF350000",x"AE000100",
x"AF360000",x"AE000100",x"AF370001",x"AE000100",x"AF370000",x"AE000100",x"AF380000",x"AE000100",
x"AF390004",x"AE000100",x"AF3A0000",x"AE000100",x"AF4803FF",x"AE000100",x"AF3D0F00",x"AE000100",
x"AF260000",x"AE000100",x"AF260800",x"AE000100",x"AF260000",x"AE000100",x"AF0B8001",x"AE000100",
x"AF0A0000",x"AE000100",x"AF0A0001",x"AE000100",x"AF0A0000",x"AE000100",x"AF260000",x"AE000100",
x"AF264000",x"AE000100",x"AF26C000",x"AE000100",x"AF264000",x"AE000100",x"AF270000",x"AE000100",
x"AF2AFE00",x"AE000100",x"AF2901FF",x"AE000100",x"AF2981FF",x"AE00FFFF",x"AF2901FF",x"AE00FFFF",
x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",
x"C0000000",x"C0010000",x"C0020000",x"C0030000",x"C0040000",x"C0050000",x"C0060000",x"C0070000",
x"C0080000",x"C0090000",x"C00A0000",x"C00B0000",x"C00C0000",x"C00D0000",x"C00E0000",x"C00F0000",
x"C0100000",x"C0110000",x"C0120000",x"C0130000",x"C0140000",x"C0150000",x"C0160000",x"C0170000",
x"C0180000",x"C0190000",x"C01A0000",x"C01B0000",x"C01C0000",x"C01D0000",x"C01E0000",x"C01F0000",
x"C0200000",x"C0210000",x"C0220000",x"C0230000",x"C0240000",x"C0250000",x"C0260000",x"C0270000",
x"C0280000",x"C0290000",x"C02A0000",x"C02B0000",x"C02C0000",x"C02D0000",x"C02E0000",x"C02F0000",
x"C0300000",x"C0310000",x"C0320000",x"C0330000",x"C0340000",x"C0350000",x"C0360000",x"C0370000",
x"C0380000",x"C0390000",x"C03A0000",x"C03B0000",x"C03C0000",x"C03D0000",x"C03E0000",x"C03F0000",
x"C0400000",x"C0410000",x"C0420000",x"C0430000",x"C0440000",x"C0450000",x"C0460000",x"C0470000",
x"C0480000",x"C0490000",x"C04A0000",x"C04B0000",x"C04C0000",x"C04D0000",x"C04E0000",x"C04F0000",
x"C0500000",x"C0510000",x"C0520000",x"C0530000",x"C0540000",x"C0550000",x"C0560000",x"C0570000",
x"C0580000",x"C0590000",x"C05A0000",x"C05B0000",x"C05C0000",x"C05D0000",x"C05E0000",x"C05F0000",
x"C0600000",x"C0610000",x"C0620000",x"C0630000",x"C0640000",x"C0650000",x"C0660000",x"C0670000",
x"C0680000",x"C0690000",x"C06A0000",x"C06B0000",x"C06C0000",x"C06D0000",x"C06E0000",x"C06F0000",
x"C0700000",x"C0710000",x"C0720000",x"C0730000",x"C0740000",x"C0750000",x"C0760000",x"C0770000",
x"C0780000",x"C0790000",x"C07A0000",x"C07B0000",x"C07C0000",x"C07D0000",x"C07E0000",x"C07F0000",
x"C0800000",x"C0810000",x"C0820000",x"C0830000",x"C0840000",x"C0850000",x"C0860000",x"C0870000",
x"C0880000",x"C0890000",x"C08A0000",x"C08B0000",x"C08C0000",x"C08D0000",x"C08E0000",x"C08F0000",
x"C0900000",x"C0910000",x"C0920000",x"C0930000",x"C0940000",x"C0950000",x"C0960000",x"C0970000",
x"C0980000",x"C0990000",x"C09A0000",x"C09B0000",x"C09C0000",x"C09D0000",x"C09E0000",x"C09F0000",
x"AF140000",x"AE000100",x"AF1E0000",x"AE000100",x"AF1F0000",x"AE000100",x"AF320000",x"AE000100",
x"AF2C0000",x"AE000100",x"AF2D0001",x"AE000100",x"AF2D0000",x"AE000100",x"AF3303FF",x"AE000100",
x"AF340000",x"AE000100",x"AF350000",x"AE000100",x"AF360003",x"AE000100",x"AF370001",x"AE000100",
x"AF370000",x"AE000100",x"AF380000",x"AE000100",x"AF390004",x"AE000100",x"AF3A0000",x"AE000100",
x"AF4803FF",x"AE000100",x"AF3D0F00",x"AE000100",x"AF260000",x"AE000100",x"AF260800",x"AE000100",
x"AF260000",x"AE000100",x"AF261080",x"AE000100",x"AF25C000",x"AE000100",x"AF4B0000",x"AE000100",
x"AF4C0003",x"AE000100",x"AF270000",x"AE000100",x"AF0B8001",x"AE000100",x"AF0A0000",x"AE000100",
x"AF0A0001",x"AE000100",x"AF0A0000",x"AE000100",x"AF3E0000",x"AE000100",x"AF460000",x"AE000100",
x"AF470000",x"AE000100",x"AF470001",x"AE000100",x"AF470000",x"AE000100",x"AF460001",x"AE000100",
x"AF27C3FF",x"AE000100",x"AF4D0450",x"AE000100",x"AF4DC450",x"AE000100",x"AF008D0E",x"AE000100",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000"
);

constant scrod_rcl_sim2_autoinit_len: integer:=81;
 
type scrod_rcl_sim2_autoinit is array (0 to scrod_rcl_sim2_autoinit_len-1) of std_logic_vector(31 downto 0);
constant init_scrod_rcl_sim2_autoinit : scrod_rcl_sim2_autoinit:=(
x"AE000010",x"AF050080",x"AE000010",x"AF060140",x"AE000010",x"AF140000",x"AE000010",x"AF1E0000",
x"AE000010",x"AF1F0000",x"AE000010",x"AF320000",x"AE000010",x"AF2C0000",x"AE000010",x"AF2D0001",
x"AE000010",x"AF2D0000",x"AE000010",x"AF3301E7",x"AE000010",x"AF340000",x"AE000010",x"AF350000",
x"AE000010",x"AF360090",x"AE000010",x"AF370001",x"AE000010",x"AF370000",x"AE000010",x"AF380020", --AF38 - lookback width at 32 windows = ~1us for sim
x"AE000010",x"AF390004",x"AE000010",x"AF3A0000",x"AE000010",x"AF4801E7",x"AE000010",x"AF3D00F0", -- default for AF3D was 0F00 but swithing to shorter ramp at 00F0
x"AE000010",x"AF260000",x"AE000010",x"AF260800",x"AE000010",x"AF260000",x"AE000010",x"AF2610E0",--x"AF2610A0", (10E0=cal mode reg - force read
x"AE000010",x"AF4B0000",x"AE000010",x"AF4C0003",x"AE000010",x"AF270000",x"AE000010",x"AF0B8001",
x"AE000010",x"AF0A0000",x"AE000010",x"AF0A0001",x"AE000010",x"AF0A0000",x"AE000010",x"AF3E0000",
x"AE000010",x"AF460000",x"AE000010",x"AF470000",x"AE000010",x"AF470001",x"AE000010",x"AF470000",
x"AE000010",x"AF460001",x"AE000010",x"AF27C1E7",x"AE000010",x"AF008D0E",x"AE000010",x"AF330002", --only readout ASIC   2
x"AF2B0FFF");-- channel mask ch 15 (0 based) should never be force readout


--x"01234567",x"AE000100",x"AF000000",x"AE000100",x"AF008000",x"AE000100",x"AE008000",x"AE000100",
--x"AE000100",x"AF00FFFF",x"AE000100",x"AE000100",x"AF008000",x"AE000100",x"AF050080",x"AE000100",
--x"AF060140",x"AE000100",
--x"AF140000",x"AE000100",x"AF1E0000",x"AE000100",x"AF1F0000",x"AE000100",x"AF320000",x"AE000100",
--x"AF2C0000",x"AE000100",x"AF2D0001",x"AE000100",x"AF2D0000",x"AE000100",x"AF3303FF",x"AE000100",
--x"AF340000",x"AE000100",x"AF350000",x"AE000100",x"AF360003",x"AE000100",x"AF370001",x"AE000100",
--x"AF370000",x"AE000100",x"AF380000",x"AE000100",x"AF390004",x"AE000100",x"AF3A0000",x"AE000100",
--x"AF4803FF",x"AE000100",x"AF3D0F00",x"AE000100",x"AF260000",x"AE000100",x"AF260800",x"AE000100",
--x"AF260000",x"AE000100",x"AF261080",x"AE000100",x"AF25C000",x"AE000100",x"AF4B0000",x"AE000100",
--x"AF4C0003",x"AE000100",x"AF270000",x"AE000100",x"AF0B8001",x"AE000100",x"AF0A0000",x"AE000100",
--x"AF0A0001",x"AE000100",x"AF0A0000",x"AE000100",x"AF3E0000",x"AE000100",x"AF460000",x"AE000100",
--x"AF470000",x"AE000100",x"AF470001",x"AE000100",x"AF470000",x"AE000100",x"AF460001",x"AE000100",
--x"AF27C3FF",x"AE000100",x"AF4D0450",x"AE000100",x"AF4DC450",x"AE000100",x"AF008D0E",x"AE000100"
--);


constant scrod_rcl_sim_autoinit_len: integer:=306;
 
type scrod_rcl_sim_autoinit is array (0 to scrod_rcl_sim_autoinit_len-1) of std_logic_vector(31 downto 0);
constant init_scrod_rcl_sim_autoinit : scrod_rcl_sim_autoinit:=(
x"01234567",x"AE000100",x"AF000000",x"AE000100",x"AF008000",x"AE000100",x"AE008000",x"AE000100",
x"AE000100",x"AF00FFFF",x"AE000100",x"AE000100",x"AF008000",x"AE000100",x"AF050080",x"AE000100",
x"AF060140",x"AE000100",x"B00005AA",x"B00205AA",x"B00405AA",x"B00605AA",x"B00805AA",x"B00A05AA",
x"AF4D0000",x"AE000100",x"AF140000",x"AE000100",x"AF1E0000",x"AE000100",x"AF320000",x"AE000100",
x"AF2C0000",x"AE000100",x"AF2D0001",x"AE000100",x"AF2D0000",x"AE000100",x"AF3303FF",x"AE000100",
x"AF340000",x"AE000100",x"AF350000",x"AE000100",x"AF360000",x"AE000100",x"AF370001",x"AE000100",
x"AF370000",x"AE000100",x"AF380000",x"AE000100",x"AF390004",x"AE000100",x"AF3A0000",x"AE000100",
x"AF4803FF",x"AE000100",x"AF3D0F00",x"AE000100",x"AF260000",x"AE000100",x"AF260800",x"AE000100",
x"AF260000",x"AE000100",x"AF0B8001",x"AE000100",x"AF0A0000",x"AE000100",x"AF0A0001",x"AE000100",
x"AF0A0000",x"AE000100",x"AF260000",x"AE000100",x"AF264000",x"AE000100",x"AF26C000",x"AE000100",
x"AF264000",x"AE000100",x"AF270000",x"AE000100",x"AF2AFE00",x"AE000100",x"AF290200",x"AE000100",
x"AF298200",x"AE00FFFF",x"AF290200",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",
x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AF4D0000",x"AE000100",x"AF140000",x"AE000100",
x"AF1E0000",x"AE000100",x"AF320000",x"AE000100",x"AF2C0000",x"AE000100",x"AF2D0001",x"AE000100",
x"AF2D0000",x"AE000100",x"AF3303FF",x"AE000100",x"AF340000",x"AE000100",x"AF350000",x"AE000100",
x"AF360000",x"AE000100",x"AF370001",x"AE000100",x"AF370000",x"AE000100",x"AF380000",x"AE000100",
x"AF390004",x"AE000100",x"AF3A0000",x"AE000100",x"AF4803FF",x"AE000100",x"AF3D0F00",x"AE000100",
x"AF260000",x"AE000100",x"AF260800",x"AE000100",x"AF260000",x"AE000100",x"AF0B8001",x"AE000100",
x"AF0A0000",x"AE000100",x"AF0A0001",x"AE000100",x"AF0A0000",x"AE000100",x"AF260000",x"AE000100",
x"AF264000",x"AE000100",x"AF26C000",x"AE000100",x"AF264000",x"AE000100",x"AF270000",x"AE000100",
x"AF2AFE00",x"AE000100",x"AF2901FF",x"AE000100",x"AF2981FF",x"AE00FFFF",x"AF2901FF",x"AE00FFFF",
x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",x"AE00FFFF",
x"AF140000",x"AE000100",x"AF1E0000",x"AE000100",x"AF1F0000",x"AE000100",x"AF320000",x"AE000100",
x"AF2C0000",x"AE000100",x"AF2D0001",x"AE000100",x"AF2D0000",x"AE000100",x"AF3303FF",x"AE000100",
x"AF340000",x"AE000100",x"AF350000",x"AE000100",x"AF360003",x"AE000100",x"AF370001",x"AE000100",
x"AF370000",x"AE000100",x"AF380000",x"AE000100",x"AF390004",x"AE000100",x"AF3A0000",x"AE000100",
x"AF4803FF",x"AE000100",x"AF3D0F00",x"AE000100",x"AF260000",x"AE000100",x"AF260800",x"AE000100",
x"AF260000",x"AE000100",x"AF261080",x"AE000100",x"AF25C000",x"AE000100",x"AF4B0000",x"AE000100",
x"AF4C0003",x"AE000100",x"AF270000",x"AE000100",x"AF0B8001",x"AE000100",x"AF0A0000",x"AE000100",
x"AF0A0001",x"AE000100",x"AF0A0000",x"AE000100",x"AF3E0000",x"AE000100",x"AF460000",x"AE000100",
x"AF470000",x"AE000100",x"AF470001",x"AE000100",x"AF470000",x"AE000100",x"AF460001",x"AE000100",
x"AF27C3FF",x"AE000100",x"AF4D0450",x"AE000100",x"AF4DC450",x"AE000100",x"AF008D0E",x"AE000100",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
x"00000000",x"00000000"
);

constant scrod_rcl_autoinit_DAC_len: integer:=181;
 
type scrod_rcl_autoinit_DAC is array (0 to scrod_rcl_autoinit_DAC_len-1) of std_logic_vector(31 downto 0);
constant init_scrod_rcl_autoinit_DAC : scrod_rcl_autoinit_DAC:=(
x"01234567",x"AE000100",x"AF000000",x"AE000100",x"AF008000",x"AE000100",x"AE008000",x"AE000100",
x"AE000100",x"AF00FFFF",x"AE000100",x"AE000100",x"AF008000",x"AE000100",x"AF050080",x"AE000100",
x"AF060140",x"AE000100",
x"C0000000",x"C0010000",x"C0020000",x"C0030000",x"C0040000",x"C0050000",x"C0060000",x"C0070000",
x"C0080000",x"C0090000",x"C00A0000",x"C00B0000",x"C00C0000",x"C00D0000",x"C00E0000",x"C00F0000",
x"C0100000",x"C0110000",x"C0120000",x"C0130000",x"C0140000",x"C0150000",x"C0160000",x"C0170000",
x"C0180000",x"C0190000",x"C01A0000",x"C01B0000",x"C01C0000",x"C01D0000",x"C01E0000",x"C01F0000",
x"C0200000",x"C0210000",x"C0220000",x"C0230000",x"C0240000",x"C0250000",x"C0260000",x"C0270000",
x"C0280000",x"C0290000",x"C02A0000",x"C02B0000",x"C02C0000",x"C02D0000",x"C02E0000",x"C02F0000",
x"C0300000",x"C0310000",x"C0320000",x"C0330000",x"C0340000",x"C0350000",x"C0360000",x"C0370000",
x"C0380000",x"C0390000",x"C03A0000",x"C03B0000",x"C03C0000",x"C03D0000",x"C03E0000",x"C03F0000",
x"C0400000",x"C0410000",x"C0420000",x"C0430000",x"C0440000",x"C0450000",x"C0460000",x"C0470000",
x"C0480000",x"C0490000",x"C04A0000",x"C04B0000",x"C04C0000",x"C04D0000",x"C04E0000",x"C04F0000",
x"C0500000",x"C0510000",x"C0520000",x"C0530000",x"C0540000",x"C0550000",x"C0560000",x"C0570000",
x"C0580000",x"C0590000",x"C05A0000",x"C05B0000",x"C05C0000",x"C05D0000",x"C05E0000",x"C05F0000",
x"C0600000",x"C0610000",x"C0620000",x"C0630000",x"C0640000",x"C0650000",x"C0660000",x"C0670000",
x"C0680000",x"C0690000",x"C06A0000",x"C06B0000",x"C06C0000",x"C06D0000",x"C06E0000",x"C06F0000",
x"C0700000",x"C0710000",x"C0720000",x"C0730000",x"C0740000",x"C0750000",x"C0760000",x"C0770000",
x"C0780000",x"C0790000",x"C07A0000",x"C07B0000",x"C07C0000",x"C07D0000",x"C07E0000",x"C07F0000",
x"C0800000",x"C0810000",x"C0820000",x"C0830000",x"C0840000",x"C0850000",x"C0860000",x"C0870000",
x"C0880000",x"C0890000",x"C08A0000",x"C08B0000",x"C08C0000",x"C08D0000",x"C08E0000",x"C08F0000",
x"C0900000",x"C0910000",x"C0920000",x"C0930000",x"C0940000",x"C0950000",x"C0960000",x"C0970000",
x"C0980000",x"C0990000",x"C09A0000",x"C09B0000",x"C09C0000",x"C09D0000",x"C09E0000",x"C09F0000",
x"AE000100",x"00000000",x"00000000"
);

 

end autoinit_definitions;

package body autoinit_definitions is

 
end autoinit_definitions;
